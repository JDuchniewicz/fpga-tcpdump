// the top module, responsible for capturing (nor now) the incoming packets
// from the network interface
module bpfcap_top(input logic clk,
                  logic reset,
                  output logic[
                  );

endmodule

